& @English:
Drills for Cannon-related 2H @English:
Cannon-related Checkmate
Red moves first and wins the game
                                                            	                   	    