 @English:
Stalemate 1G @English:
Flanking Trio Checkmate
Red moves first and wins the game
                                        
                      	     
	      		        