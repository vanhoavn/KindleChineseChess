 @English:
Horse – Cannon 3J @English:
Horse – Cannon Checkmate
Red moves first and wins the game
                                                                 	      	                