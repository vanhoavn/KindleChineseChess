 @English:
Chariot and Pawn 5J @English:
Chariot and Pawn Checkmate
Red moves first and wins the game
                                                                     	             	          	   		        