' @English:
Drills for Chariot Related 2I @English:
Chariot Related Checkmate
Red moves first and wins the game
                                                             
                   	      