' @English:
Chariot and Double Cannons 6T @English:
Chariot and Double Cannons Checkmate
Red moves first and wins the game
                                                              	    
	  
       			  