 @English:
Angler Horse 2F @English:
Angler Horse Checkmate
Red moves first and wins the game
                                                        
       	    
	         