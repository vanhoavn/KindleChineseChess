+ @English:
Double Devils Knocking at Door 1Z @English:
"Double Devils Knocking at Door" Checkmate
Red moves first and wins the game
                                                         
       	      
 	   	       