 @English:
Chariot and Cannon 4L @English:
Chariot and Cannon Checkmate
Red moves first and wins the game
                                       
                  		                             