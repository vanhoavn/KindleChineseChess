 @English:
Flanking Trio 3G @English:
Flanking Trio Checkmate
Red moves first and wins the game
                                        
                      	     
	      		        