1 @English:
Drills for Horse and Cannon Combined 7S @English:
Horse and Cannon Combined Checkmate
Red moves first and wins the game
                                                                         		                   