% @English:
Chariot, Cannon and Pawn 2R @English:
Chariot, Cannon and Pawn Checkmate
Red moves first and wins the game
                                                                        
                   