 @English:
Horse and Cannon 2J @English:
Horse and Cannon Checkmate
Red moves first and wins the game
                                                                           
  
         