' @English:
Drills for Chariot Related 8I @English:
Chariot Related Checkmate
Red moves first and wins the game
                                                                                          