 @English:
Palcorner Horse 3I @English:
Palcorner Horse Checkmate
Red moves first and wins the game
                                                              
   	     
    	       