# @English:
Chariot-Horse Zugzwang 4k @English:
Chariot-Horse Zugzwang Checkmate (White Horse Showing Hoof)
Red moves first and wins the game
                                                      
        	      	 
  			        