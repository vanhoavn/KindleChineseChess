$ @English:
Chariot, Horse and Pawn 7Q @English:
Chariot, Horse and Pawn Checkmate
Red moves first and wins the game
                                      
               
       	        	         