 @English:
Iron-Bolt 2C @English:
Iron-Bolt Checkmate
Red moves first and wins the game
                                                   
           	      	
  			      