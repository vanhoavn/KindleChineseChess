 @English:
Double Cannon 1G @English:
Double Cannon Checkmate
Red moves first and wins the game
                                                         
        	     
	   	           