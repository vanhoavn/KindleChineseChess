4 @English:
Drills for Chariot and Cannon Combined 16U @English:
Chariot and Cannon Combined Checkmate
Red moves first and wins the game
                                                                        		      	   