 @English:
Horse – Cannon 2J @English:
Horse – Cannon Checkmate
Red moves first and wins the game
                                                      
             
    	        