* @English:
Drills for Chariot and Horse 15K @English:
Chariot and Horse Checkmate
Red moves first and wins the game
                                                           
             		       	 