+ @English:
Double Devils Knocking at Door 2Z @English:
"Double Devils Knocking at Door" Checkmate
Red moves first and wins the game
                                                                                  		   