& @English:
Chariot, Horse and Cannon 4S @English:
Chariot, Horse and Cannon Checkmate
Red moves first and wins the game
                                                               	     
	 
    