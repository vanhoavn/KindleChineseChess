, @English:
Chariot, Horse, Cannon and Pawn 2Y @English:
Chariot, Horse, Cannon and Pawn Checkmate
Red moves first and wins the game
                                                         	             	          