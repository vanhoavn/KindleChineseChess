+ @English:
Chariot-Horse (BA-Huang Horse) 1X @English:
Chariot-Horse (BA-Huang Horse) Checkmate
Red moves first and wins the game
                                                         
       	     
	            