$ @English:
Chariot-Cannon Discover 1Q @English:
Chariot-Cannon Discover Checkmate
Red moves first and wins the game
                                                                       		                  