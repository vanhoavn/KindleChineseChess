 @English:
Smothered 1C @English:
Smothered Checkmate
Red moves first and wins the game
                                                                                    