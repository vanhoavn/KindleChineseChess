 @English:
Smothered 3C @English:
Smothered Checkmate
Red moves first and wins the game
                                                                      
		
  	       