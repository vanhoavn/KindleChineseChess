& @English:
Chariot, Horse and Cannon 2S @English:
Chariot, Horse and Cannon Checkmate
Red moves first and wins the game
                                                          
             
	        