& @English:
Drills for Cannon-related 3H @English:
Cannon-related Checkmate
Red moves first and wins the game
                                                                                       