 @English:
Horse-Pawn 1D @English:
Horse-Pawn Checkmate
Red moves first and wins the game
                                                                                     	 