& @English:
Drills for Cannon-related 1H @English:
Cannon-related Checkmate
Red moves first and wins the game
                                                                                