$ @English:
Chariot, Horse and Pawn 3Q @English:
Chariot, Horse and Pawn Checkmate
Red moves first and wins the game
                                                       	
       	         
              