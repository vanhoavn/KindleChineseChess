# @English:
Horse, Cannon and Pawn 8P @English:
Horse, Cannon and Pawn Checkmate
Red moves first and wins the game
                                                      
                                