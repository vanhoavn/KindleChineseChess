# @English:
Horse, Cannon and Pawn 2P @English:
Horse, Cannon and Pawn Checkmate
Red moves first and wins the game
                                                         	
	                  