% @English:
Chariot, Cannon and Pawn 3R @English:
Chariot, Cannon and Pawn Checkmate
Red moves first and wins the game
                                                                  	             		   