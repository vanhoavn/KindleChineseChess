 @English:
Cannon-Pawn 1E @English:
Cannon-Pawn Checkmate
Red moves first and wins the game
                                                                    	      	    			   		  		 