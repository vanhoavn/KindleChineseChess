 @English:
Double Horses 2G @English:
Double Horses Checkmate
Red moves first and wins the game
                                                                           	 
             