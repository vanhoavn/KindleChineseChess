 @English:
Octagonal Horse 2I @English:
Octagonal Horse Checkmate
Red moves first and wins the game
                                                                                   						     