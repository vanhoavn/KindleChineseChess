 @English:
Double Chariots 5I @English:
Double Chariots Checkmate
Red moves first and wins the game
                                        
                 	
            	      	     	  