" @English:
Face-to-Face Laughing 3O @English:
Face-to-Face Laughing Checkmate
Red moves first and wins the game
                                                                     	              		 