" @English:
Face-to-Face Laughing 1O @English:
Face-to-Face Laughing Checkmate
Red moves first and wins the game
                                                                           
 	
    