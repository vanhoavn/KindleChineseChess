 @English:
Double Cannons 4H @English:
Double Cannons Checkmate
Red moves first and wins the game
                                                                                         