 @English:
Cannon-Pawn 5E @English:
Cannon-Pawn Checkmate
Red moves first and wins the game
                                                                             
 	        	 		   	 		  	 	 	  	 	   