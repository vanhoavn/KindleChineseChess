 @English:
Cannon-Pawn 4E @English:
Cannon-Pawn Checkmate
Red moves first and wins the game
                                                                                  		 	     	    		 