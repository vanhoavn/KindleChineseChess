 @English:
Chariot and Cannon 3L @English:
Chariot and Cannon Checkmate
Red moves first and wins the game
                                                                  	      	
  		       	     