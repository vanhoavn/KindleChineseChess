 @English:
Horse-Pawn 3D @English:
Horse-Pawn Checkmate
Red moves first and wins the game
                                                                        
   
      		 	                          