 @English:
Chariot and Cannon 1L @English:
Chariot and Cannon Checkmate
Red moves first and wins the game
                                                                 	        	         