% @English:
Drills for Horse-Related 7G @English:
Horse-Related Checkmate
Red moves first and wins the game
                                                                   	         
      