 @English:
Horse-Pawn 4D @English:
Horse-Pawn Checkmate
Red moves first and wins the game
                                                                                        