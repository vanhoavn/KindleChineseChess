 @English:
Cannon Smothered 2J @English:
Cannon Smothered Checkmate
Red moves first and wins the game
                                                                  	           	       