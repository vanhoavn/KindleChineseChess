  @English:
Simultaneous Double 3M @English:
Simultaneous Double Checkmate
Red moves first and wins the game
                                                                       		     