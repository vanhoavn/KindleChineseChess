 @English:
Throat-cutting 3H @English:
Throat-cutting Checkmate
Red moves first and wins the game
                                                                	            	        