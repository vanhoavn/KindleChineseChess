 @English:
Horse and Cannon 8J @English:
Horse and Cannon Checkmate
Red moves first and wins the game
                                                            	        	        
  						 