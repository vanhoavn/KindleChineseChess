& @English:
Chariot, Horse and Cannon 8S @English:
Chariot, Horse and Cannon Checkmate
Red moves first and wins the game
                                                                 	       	
                     	 