' @English:
Drills for Chariot Related 1I @English:
Chariot Related Checkmate
Red moves first and wins the game
                                         
             
  	                	  	     