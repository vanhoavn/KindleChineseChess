 @English:
Double Chariots 3I @English:
Double Chariots Checkmate
Red moves first and wins the game
                                                      
        	      
	             