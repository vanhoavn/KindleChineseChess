 @English:
Horse and Cannon 3J @English:
Horse and Cannon Checkmate
Red moves first and wins the game
                                                                                      