 @English:
Double Chariots 1I @English:
Double Chariots Checkmate
Red moves first and wins the game
                                                                   	       	                  