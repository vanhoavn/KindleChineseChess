% @English:
Double Chariots and Pawn 2R @English:
Double Chariots and Pawn Checkmate
Red moves first and wins the game
                                                                        
		
 		         