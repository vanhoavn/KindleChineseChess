& @English:
Chariot and Double Horses 5S @English:
Chariot and Double Horses Checkmate
Red moves first and wins the game
                                                          	  
    	                	     