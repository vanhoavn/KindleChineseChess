 @English:
Throat-cutting 1H @English:
Throat-cutting Checkmate
Red moves first and wins the game
                                                                 	           	    	      