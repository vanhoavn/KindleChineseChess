$ @English:
Double Cannons and Pawn 3Q @English:
Double Cannons and Pawn Checkmate
Red moves first and wins the game
                                                         
        	    
	   			 	  