% @English:
Chariot, Cannon and Pawn 7R @English:
Chariot, Cannon and Pawn Checkmate
Red moves first and wins the game
                                                          	            
                   