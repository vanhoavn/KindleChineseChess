 @English:
Horse-Pawn 5D @English:
Horse-Pawn Checkmate
Red moves first and wins the game
                                                                                              