 @English:
Double Cannon 2G @English:
Double Cannon Checkmate
Red moves first and wins the game
                                                               	      
	 
      