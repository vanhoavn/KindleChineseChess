 @English:
Exposed Cannon 1H @English:
Exposed Cannon Checkmate
Red moves first and wins the game
                                                         
    	     
	        