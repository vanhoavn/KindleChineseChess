& @English:
Chariot and Double Horses 6S @English:
Chariot and Double Horses Checkmate
Red moves first and wins the game
                                        
                              
		            