 @English:
Chariot and Pawn 4J @English:
Chariot and Pawn Checkmate
Red moves first and wins the game
                                                             
                    	          