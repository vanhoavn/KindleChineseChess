A @English:
Drills for Chariot, Cannon, Horse and Pawn Combined 12b @English:
Chariot, Cannon, Horse and Pawn Combined Checkmate
Red moves first and wins the game
                                                             	       	           