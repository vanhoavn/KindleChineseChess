' @English:
Chariot and Double Cannons 2T @English:
Chariot and Double Cannons Checkmate
Red moves first and wins the game
                                                                	     
	 
              	  