% @English:
Chariot, Cannon and Pawn 6R @English:
Chariot, Cannon and Pawn Checkmate
Red moves first and wins the game
                                                           
     	     
	     	              