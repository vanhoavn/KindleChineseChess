' @English:
Chariot and Double Cannons 5T @English:
Chariot and Double Cannons Checkmate
Red moves first and wins the game
                                                             
                     	          