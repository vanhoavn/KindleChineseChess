$ @English:
Double Cannons and Pawn 4Q @English:
Double Cannons and Pawn Checkmate
Red moves first and wins the game
                                                        
                          