 @English:
Tiger Silhouette 3J @English:
Tiger Silhouette Checkmate
Red moves first and wins the game
                                           
              
      	        	         			  