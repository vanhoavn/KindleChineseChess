& @English:
Drills for Cannon-related 6H @English:
Cannon-related Checkmate
Red moves first and wins the game
                                       
                  
                   