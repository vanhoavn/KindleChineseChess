% @English:
Drills for Horse-Related 5G @English:
Horse-Related Checkmate
Red moves first and wins the game
                                                                                        