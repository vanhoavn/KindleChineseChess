& @English:
Chariot, Horse and Cannon 9S @English:
Chariot, Horse and Cannon Checkmate
Red moves first and wins the game
                                                         
      	        	             