1 @English:
Drills for Horse and Cannon Combined 9S @English:
Horse and Cannon Combined Checkmate
Red moves first and wins the game
                                                                                                  