 @English:
Chariot and Pawn 3J @English:
Chariot and Pawn Checkmate
Red moves first and wins the game
                                                            
       	     	   		    