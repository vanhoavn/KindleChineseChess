 @English:
Palcorner Horse 1I @English:
Palcorner Horse Checkmate
Red moves first and wins the game
                                                         
        	   
	        