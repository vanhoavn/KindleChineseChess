 @English:
Elbow Horse 1E @English:
Elbow Horse Checkmate
Red moves first and wins the game
                                                                             	 