 @English:
Elbow Horse 3E @English:
Elbow Horse Checkmate
Red moves first and wins the game
                                        
               
                         