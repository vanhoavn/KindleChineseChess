 @English:
Tiger Silhouette 1J @English:
Tiger Silhouette Checkmate
Red moves first and wins the game
                                                         
       	     
	        	       