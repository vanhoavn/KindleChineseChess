 @English:
Elbow Horse 2E @English:
Elbow Horse Checkmate
Red moves first and wins the game
                                                                              			      