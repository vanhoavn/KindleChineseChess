% @English:
Double Chariots and Pawn 3R @English:
Double Chariots and Pawn Checkmate
Red moves first and wins the game
                                                                      
              