 @English:
Double Cannons 1H @English:
Double Cannons Checkmate
Red moves first and wins the game
                                                                           
  
      	 	  