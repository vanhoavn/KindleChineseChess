 @English:
Horse – Cannon 1J @English:
Horse – Cannon Checkmate
Red moves first and wins the game
                                                           	 	                        