' @English:
Drills for Chariot Related 4I @English:
Chariot Related Checkmate
Red moves first and wins the game
                                                            
              
        