 @English:
Double Horses 4G @English:
Double Horses Checkmate
Red moves first and wins the game
                                                                  	       	                 