& @English:
Drills for Cannon-related 8H @English:
Cannon-related Checkmate
Red moves first and wins the game
                                                                                            