 @English:
Horse and Cannon 4J @English:
Horse and Cannon Checkmate
Red moves first and wins the game
                                                                        
		                