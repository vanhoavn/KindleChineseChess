& @English:
Drills for Cannon-related 4H @English:
Cannon-related Checkmate
Red moves first and wins the game
                                                             	                     		   		 