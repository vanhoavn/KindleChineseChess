$ @English:
Chariot-Cannon Discover 2Q @English:
Chariot-Cannon Discover Checkmate
Red moves first and wins the game
                                                      
        	       	
                  