 @English:
Double Cannons 2H @English:
Double Cannons Checkmate
Red moves first and wins the game
                                                           
       	      
      		   	   