) @English:
Heavenly and Earthly Cannons 3V @English:
Heavenly and Earthly Cannons Checkmate
Red moves first and wins the game
                                                                     
		             		    