% @English:
Drills for Horse-Related 8G @English:
Horse-Related Checkmate
Red moves first and wins the game
                                          
                     
                   			 	 