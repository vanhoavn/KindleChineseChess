 @English:
Double Cannon 3G @English:
Double Cannon Checkmate
Red moves first and wins the game
                                                      	
	              
         