 @English:
Double Horses 5G @English:
Double Horses Checkmate
Red moves first and wins the game
                                                              
            		
    								  