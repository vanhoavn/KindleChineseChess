# @English:
Double Horses and Pawn 5P @English:
Double Horses and Pawn Checkmate
Red moves first and wins the game
                                                                                				 