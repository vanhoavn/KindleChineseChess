% @English:
Drills for Horse-Related 4G @English:
Horse-Related Checkmate
Red moves first and wins the game
                                                                               	      