 @English:
Octagonal Horse 1I @English:
Octagonal Horse Checkmate
Red moves first and wins the game
                                                                   	       	            