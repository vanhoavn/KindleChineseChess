% @English:
Drills for Horse-Related 3G @English:
Horse-Related Checkmate
Red moves first and wins the game
                                                                                 	  