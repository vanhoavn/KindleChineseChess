 @English:
Chariot and Pawn 2J @English:
Chariot and Pawn Checkmate
Red moves first and wins the game
                                                                                  !        				  	               