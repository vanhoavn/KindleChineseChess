  @English:
Simultaneous Double 1M @English:
Simultaneous Double Checkmate
Red moves first and wins the game
                                                                                