# @English:
Double Horses and Pawn 4P @English:
Double Horses and Pawn Checkmate
Red moves first and wins the game
                                    
               
    	                   	 	   	 