' @English:
Drills for Chariot Related 6I @English:
Chariot Related Checkmate
Red moves first and wins the game
                                                                                         