" @English:
Face-to-Face Laughing 4O @English:
Face-to-Face Laughing Checkmate
Red moves first and wins the game
                                                                               	 	  