) @English:
Drills for Chariot and Horse 2K @English:
Chariot and Horse Checkmate
Red moves first and wins the game
                                                             	       	           	    