# @English:
Double Horses and Pawn 2P @English:
Double Horses and Pawn Checkmate
Red moves first and wins the game
                                                                    	       	        