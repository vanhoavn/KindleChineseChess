' @English:
Drills for Chariot Related 3I @English:
Chariot Related Checkmate
Red moves first and wins the game
                                                          		                              