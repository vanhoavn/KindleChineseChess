 @English:
Double Horses 1G @English:
Double Horses Checkmate
Red moves first and wins the game
                                           
              
        	      	         