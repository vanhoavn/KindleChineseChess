 @English:
Iron-Bolt 1C @English:
Iron-Bolt Checkmate
Red moves first and wins the game
                                                          
        	       	
    	  