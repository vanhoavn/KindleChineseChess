 @English:
Cannon Smothered 4J @English:
Cannon Smothered Checkmate
Red moves first and wins the game
                                                                       	    	    	   	     