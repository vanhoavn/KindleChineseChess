 @English:
Stalemate 2C @English:
Stalemate Checkmate
Red moves first and wins the game
                                                                                   	   	   