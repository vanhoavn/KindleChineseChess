# @English:
Repatriation of Buddha 2P @English:
Repatriation of Buddha Checkmate
Red moves first and wins the game
                                                       
             
	              