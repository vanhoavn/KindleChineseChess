 @English:
Double Cannons 3H @English:
Double Cannons Checkmate
Red moves first and wins the game
                                       
                                        	 