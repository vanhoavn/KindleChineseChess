' @English:
Drills for Chariot Related 7I @English:
Chariot Related Checkmate
Red moves first and wins the game
                                                         
 
                               