" @English:
Face-to-Face Laughing 2O @English:
Face-to-Face Laughing Checkmate
Red moves first and wins the game
                                                                     
		
          