% @English:
Drills for Horse-Related 6G @English:
Horse-Related Checkmate
Red moves first and wins the game
                                                         
                          