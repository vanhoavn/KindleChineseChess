& @English:
Drills for Cannon-related 5H @English:
Cannon-related Checkmate
Red moves first and wins the game
                                                              	                     	  