 @English:
Flanking Trio 2G @English:
Flanking Trio Checkmate
Red moves first and wins the game
                                      
                          	    
	                