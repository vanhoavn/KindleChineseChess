4 @English:
Drills for Chariot and Cannon Combined 15U @English:
Chariot and Cannon Combined Checkmate
Red moves first and wins the game
                                                       
	               	
 		       		    