 @English:
Cannon-Pawn 3E @English:
Cannon-Pawn Checkmate
Red moves first and wins the game
                                                                                   						 	 