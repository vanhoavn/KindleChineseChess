 @English:
Cannon-Pawn 2E @English:
Cannon-Pawn Checkmate
Red moves first and wins the game
                                            
              	                                			 