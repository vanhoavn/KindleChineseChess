 @English:
Double Horses 3G @English:
Double Horses Checkmate
Red moves first and wins the game
                                                        	 	                           