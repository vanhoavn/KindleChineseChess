 @English:
Palcorner Horse 2I @English:
Palcorner Horse Checkmate
Red moves first and wins the game
                                                                	     
	   	        		     	 