 @English:
Angler Horse 3F @English:
Angler Horse Checkmate
Red moves first and wins the game
                                                     
    	  
          	           		     