 @English:
Angler Horse 1F @English:
Angler Horse Checkmate
Red moves first and wins the game
                                                                  	     
 	
               