 @English:
Smothered 2C @English:
Smothered Checkmate
Red moves first and wins the game
                                                                    	        	    