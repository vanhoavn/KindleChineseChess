# @English:
Chariot-Horse Zugzwang 1k @English:
Chariot-Horse Zugzwang Checkmate (White Horse Showing Hoof)
Red moves first and wins the game
                                                          
        	    	 
  	           