 @English:
Chariot and Cannon 2L @English:
Chariot and Cannon Checkmate
Red moves first and wins the game
                                                           
      	     
	         		    