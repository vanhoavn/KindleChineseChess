 @English:
Horse and Cannon 5J @English:
Horse and Cannon Checkmate
Red moves first and wins the game
                                                                                    ! 		 	 	      