 @English:
Double Cannons 5H @English:
Double Cannons Checkmate
Red moves first and wins the game
                                                                    	            		                       