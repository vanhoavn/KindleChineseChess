 @English:
Octagonal Horse 3I @English:
Octagonal Horse Checkmate
Red moves first and wins the game
                                                             
  
               	    