) @English:
Drills for Chariot and Horse 9K @English:
Chariot and Horse Checkmate
Red moves first and wins the game
                                                         
              	 
  	       