& @English:
Drills for Cannon-related 7H @English:
Cannon-related Checkmate
Red moves first and wins the game
                                                                	               