 @English:
Cannon Smothered 1J @English:
Cannon Smothered Checkmate
Red moves first and wins the game
                                       
   
              	       	                   