# @English:
Repatriation of Buddha 3P @English:
Repatriation of Buddha Checkmate
Red moves first and wins the game
                                                    
        	        	
       