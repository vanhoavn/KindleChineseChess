 @English:
Throat-cutting 2H @English:
Throat-cutting Checkmate
Red moves first and wins the game
                                                                        
		                     