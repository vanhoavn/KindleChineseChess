 @English:
Double Chariots 2I @English:
Double Chariots Checkmate
Red moves first and wins the game
                                                             
       	    	      	      