 @English:
Double Chariots 4I @English:
Double Chariots Checkmate
Red moves first and wins the game
                                                       
                    
                  		   