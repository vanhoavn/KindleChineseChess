@ @English:
Drills for Chariot, Cannon, Horse and Pawn Combined 3b @English:
Chariot, Cannon, Horse and Pawn Combined Checkmate
Red moves first and wins the game
                                                          	     	                 