$ @English:
Chariot-Cannon Discover 3Q @English:
Chariot-Cannon Discover Checkmate
Red moves first and wins the game
                                      
                           
		                            