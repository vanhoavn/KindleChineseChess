 @English:
Horse-Pawn 6D @English:
Horse-Pawn Checkmate
Red moves first and wins the game
                                                                    	       	            