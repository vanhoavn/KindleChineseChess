# @English:
Horse, Cannon and Pawn 9P @English:
Horse, Cannon and Pawn Checkmate
Red moves first and wins the game
                                                                  	       	          				 