' @English:
Chariot and Double Cannons 3T @English:
Chariot and Double Cannons Checkmate
Red moves first and wins the game
                                                            
   	        	
 %   	   	               