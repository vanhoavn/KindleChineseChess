3 @English:
Drills for Chariot and Cannon Combined 5U @English:
Chariot and Cannon Combined Checkmate
Red moves first and wins the game
                                                         
             
               