 @English:
Chariot and Pawn 1J @English:
Chariot and Pawn Checkmate
Red moves first and wins the game
                                                              
      	             