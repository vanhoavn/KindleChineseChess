$ @English:
Chariot, Horse and Pawn 4Q @English:
Chariot, Horse and Pawn Checkmate
Red moves first and wins the game
                                         
                         	      	
 	  	     		 