 @English:
Horse and Cannon 6J @English:
Horse and Cannon Checkmate
Red moves first and wins the game
                                                                  
          
  		      