$ @English:
Chariot, Horse and Pawn 8Q @English:
Chariot, Horse and Pawn Checkmate
Red moves first and wins the game
                                                        	             
	 
    	        		 