 @English:
Stalemate 3C @English:
Stalemate Checkmate
Red moves first and wins the game
                                                            
                  
    	 		 