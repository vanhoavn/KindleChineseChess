) @English:
Heavenly and Earthly Cannons 2V @English:
Heavenly and Earthly Cannons Checkmate
Red moves first and wins the game
                                                        
       	     
	     				  	     