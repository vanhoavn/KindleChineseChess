@ @English:
Drills for Chariot, Cannon, Horse and Pawn Combined 6b @English:
Chariot, Cannon, Horse and Pawn Combined Checkmate
Red moves first and wins the game
                                                      
       	     	   	    		   