% @English:
Drills for Horse-Related 1G @English:
Horse-Related Checkmate
Red moves first and wins the game
                                             
               	              	     