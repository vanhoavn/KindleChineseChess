  @English:
Simultaneous Double 2M @English:
Simultaneous Double Checkmate
Red moves first and wins the game
                                                                                  