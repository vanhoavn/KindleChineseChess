- @English:
Chariot, Horse, Cannon and Pawn 10Y @English:
Chariot, Horse, Cannon and Pawn Checkmate
Red moves first and wins the game
                                                               	   
	    	        