' @English:
Drills for Chariot Related 5I @English:
Chariot Related Checkmate
Red moves first and wins the game
                                                                         
	        