 @English:
Chariot and Cannon 5L @English:
Chariot and Cannon Checkmate
Red moves first and wins the game
                                                               	                       		 							 