 @English:
Horse and Cannon 7J @English:
Horse and Cannon Checkmate
Red moves first and wins the game
                                                           	           
      !  			 		   		     	 