, @English:
Fishing the Moon Under Deep Sea 2Y @English:
Fishing-the-Moon-Under-Deep-Sea Checkmate
Red moves first and wins the game
                                                            	                                        