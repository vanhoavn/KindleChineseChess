 @English:
Tiger Silhouette 2J @English:
Tiger Silhouette Checkmate
Red moves first and wins the game
                                                         
      	      
	   	            