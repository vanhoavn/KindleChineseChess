 @English:
Cannon Smothered 3J @English:
Cannon Smothered Checkmate
Red moves first and wins the game
                                          
                           	       	  