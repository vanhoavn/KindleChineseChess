& @English:
Chariot and Double Horses 2S @English:
Chariot and Double Horses Checkmate
Red moves first and wins the game
                                        
                 	
               	             