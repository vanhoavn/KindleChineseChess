# @English:
Repatriation of Buddha 1P @English:
Repatriation of Buddha Checkmate
Red moves first and wins the game
                                                                    	      	              