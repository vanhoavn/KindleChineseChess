 @English:
Exposed Cannon 2H @English:
Exposed Cannon Checkmate
Red moves first and wins the game
                                                        
       	      	       