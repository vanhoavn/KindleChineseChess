$ @English:
Double Cannons and Pawn 2Q @English:
Double Cannons and Pawn Checkmate
Red moves first and wins the game
                                                           
                         