% @English:
Double Chariots and Pawn 4R @English:
Double Chariots and Pawn Checkmate
Red moves first and wins the game
                                                       
      	        	             		 