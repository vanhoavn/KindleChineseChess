 @English:
Iron-Bolt 3C @English:
Iron-Bolt Checkmate
Red moves first and wins the game
                                                                                     		   