 @English:
Chariot and Cannon 6L @English:
Chariot and Cannon Checkmate
Red moves first and wins the game
                                                                    	     
      	  