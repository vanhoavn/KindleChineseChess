 @English:
Horse-Pawn 2D @English:
Horse-Pawn Checkmate
Red moves first and wins the game
                                                                       
   
  	 		 				 