% @English:
Drills for Horse-Related 2G @English:
Horse-Related Checkmate
Red moves first and wins the game
                                                                                     	      