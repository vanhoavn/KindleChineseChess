 @English:
Horse and Cannon 1J @English:
Horse and Cannon Checkmate
Red moves first and wins the game
                                                              	               	    